/*
	this file is included by index.cgi
*/


var TITLE = «zasm - z80 assembler - download page»

var DESCRIPTION =
«zasm - z80 assembler - zasm is a command line z80 assembler for unix-style operating systems.
it is available as source and some precompiled binaries, e.g. for Linux and MacOS X.
it creates output in binary or intel hex file format and can create
some special formats for ZX Spectrum emulators, e.g. ".TAP" and ".SNA" files.»

var KEYWORDS = «zasm, z80 assembler, ZX Spectrum, kio»

var ROBOTS = «index,follow»


var MAIN = 
«
h4	Source of 'zasm' - z80 assembler
p.center Documentation is in <a href="Documentation/">Documentation/</a> and tarballs are in <a href="Distributions/">Distributions/</a>.
		Source can also be checked out from <a href="/Git/">the Git</a>.
		A cgi interface for online assembling is at <a href="/cgi-bin/zasm.cgi">/cgi-bin/zasm.cgi</a>.
»


